module TransRecLogic_tb ();
reg [7:0] TxDat;
reg pclk, clr_b, t_empty, r_full;    
wire [7:0] RxData;
wire read_en, inc_ptr;


    
    
endmodule

