module alu(
    input
    output
)