module cpu_top (
    input reset,
    input disable_cpu_clock,
    input clock,
    input clr_mem,
)

endmodule